module CarryWaveGen (
  input clk,
  input rst,
  output reg [9:0] SinWave,
  output reg [9:0] CosWave
  );

  reg [7:0] count=0;

  always @ ( posedge clk or posedge rst ) begin
    if (rst) begin
      count = 0;
    end else begin
      if (count == 199) begin
        count = 0;
      end else begin
        count = count + 1;
      end
    end

    case (count)
    0:begin SinWave<=0;CosWave<=399; end
    1:begin SinWave<=13;CosWave<=399; end
    2:begin SinWave<=25;CosWave<=398; end
    3:begin SinWave<=38;CosWave<=397; end
    4:begin SinWave<=50;CosWave<=396; end
    5:begin SinWave<=62;CosWave<=394; end
    6:begin SinWave<=75;CosWave<=392; end
    7:begin SinWave<=87;CosWave<=389; end
    8:begin SinWave<=99;CosWave<=386; end
    9:begin SinWave<=111;CosWave<=383; end
    10:begin SinWave<=123;CosWave<=379; end
    11:begin SinWave<=135;CosWave<=375; end
    12:begin SinWave<=147;CosWave<=371; end
    13:begin SinWave<=158;CosWave<=366; end
    14:begin SinWave<=170;CosWave<=361; end
    15:begin SinWave<=181;CosWave<=356; end
    16:begin SinWave<=192;CosWave<=350; end
    17:begin SinWave<=203;CosWave<=343; end
    18:begin SinWave<=214;CosWave<=337; end
    19:begin SinWave<=224;CosWave<=330; end
    20:begin SinWave<=235;CosWave<=323; end
    21:begin SinWave<=245;CosWave<=315; end
    22:begin SinWave<=254;CosWave<=307; end
    23:begin SinWave<=264;CosWave<=299; end
    24:begin SinWave<=273;CosWave<=291; end
    25:begin SinWave<=282;CosWave<=282; end
    26:begin SinWave<=291;CosWave<=273; end
    27:begin SinWave<=299;CosWave<=264; end
    28:begin SinWave<=307;CosWave<=254; end
    29:begin SinWave<=315;CosWave<=245; end
    30:begin SinWave<=323;CosWave<=235; end
    31:begin SinWave<=330;CosWave<=224; end
    32:begin SinWave<=337;CosWave<=214; end
    33:begin SinWave<=343;CosWave<=203; end
    34:begin SinWave<=350;CosWave<=192; end
    35:begin SinWave<=356;CosWave<=181; end
    36:begin SinWave<=361;CosWave<=170; end
    37:begin SinWave<=366;CosWave<=158; end
    38:begin SinWave<=371;CosWave<=147; end
    39:begin SinWave<=375;CosWave<=135; end
    40:begin SinWave<=379;CosWave<=123; end
    41:begin SinWave<=383;CosWave<=111; end
    42:begin SinWave<=386;CosWave<=99; end
    43:begin SinWave<=389;CosWave<=87; end
    44:begin SinWave<=392;CosWave<=75; end
    45:begin SinWave<=394;CosWave<=62; end
    46:begin SinWave<=396;CosWave<=50; end
    47:begin SinWave<=397;CosWave<=38; end
    48:begin SinWave<=398;CosWave<=25; end
    49:begin SinWave<=399;CosWave<=13; end
    50:begin SinWave<=399;CosWave<=0; end
    51:begin SinWave<=399;CosWave<=-13; end
    52:begin SinWave<=398;CosWave<=-25; end
    53:begin SinWave<=397;CosWave<=-38; end
    54:begin SinWave<=396;CosWave<=-50; end
    55:begin SinWave<=394;CosWave<=-62; end
    56:begin SinWave<=392;CosWave<=-75; end
    57:begin SinWave<=389;CosWave<=-87; end
    58:begin SinWave<=386;CosWave<=-99; end
    59:begin SinWave<=383;CosWave<=-111; end
    60:begin SinWave<=379;CosWave<=-123; end
    61:begin SinWave<=375;CosWave<=-135; end
    62:begin SinWave<=371;CosWave<=-147; end
    63:begin SinWave<=366;CosWave<=-158; end
    64:begin SinWave<=361;CosWave<=-170; end
    65:begin SinWave<=356;CosWave<=-181; end
    66:begin SinWave<=350;CosWave<=-192; end
    67:begin SinWave<=343;CosWave<=-203; end
    68:begin SinWave<=337;CosWave<=-214; end
    69:begin SinWave<=330;CosWave<=-224; end
    70:begin SinWave<=323;CosWave<=-235; end
    71:begin SinWave<=315;CosWave<=-245; end
    72:begin SinWave<=307;CosWave<=-254; end
    73:begin SinWave<=299;CosWave<=-264; end
    74:begin SinWave<=291;CosWave<=-273; end
    75:begin SinWave<=282;CosWave<=-282; end
    76:begin SinWave<=273;CosWave<=-291; end
    77:begin SinWave<=264;CosWave<=-299; end
    78:begin SinWave<=254;CosWave<=-307; end
    79:begin SinWave<=245;CosWave<=-315; end
    80:begin SinWave<=235;CosWave<=-323; end
    81:begin SinWave<=224;CosWave<=-330; end
    82:begin SinWave<=214;CosWave<=-337; end
    83:begin SinWave<=203;CosWave<=-343; end
    84:begin SinWave<=192;CosWave<=-350; end
    85:begin SinWave<=181;CosWave<=-356; end
    86:begin SinWave<=170;CosWave<=-361; end
    87:begin SinWave<=158;CosWave<=-366; end
    88:begin SinWave<=147;CosWave<=-371; end
    89:begin SinWave<=135;CosWave<=-375; end
    90:begin SinWave<=123;CosWave<=-379; end
    91:begin SinWave<=111;CosWave<=-383; end
    92:begin SinWave<=99;CosWave<=-386; end
    93:begin SinWave<=87;CosWave<=-389; end
    94:begin SinWave<=75;CosWave<=-392; end
    95:begin SinWave<=62;CosWave<=-394; end
    96:begin SinWave<=50;CosWave<=-396; end
    97:begin SinWave<=38;CosWave<=-397; end
    98:begin SinWave<=25;CosWave<=-398; end
    99:begin SinWave<=13;CosWave<=-399; end
    100:begin SinWave<=0;CosWave<=-399; end
    101:begin SinWave<=-13;CosWave<=-399; end
    102:begin SinWave<=-25;CosWave<=-398; end
    103:begin SinWave<=-38;CosWave<=-397; end
    104:begin SinWave<=-50;CosWave<=-396; end
    105:begin SinWave<=-62;CosWave<=-394; end
    106:begin SinWave<=-75;CosWave<=-392; end
    107:begin SinWave<=-87;CosWave<=-389; end
    108:begin SinWave<=-99;CosWave<=-386; end
    109:begin SinWave<=-111;CosWave<=-383; end
    110:begin SinWave<=-123;CosWave<=-379; end
    111:begin SinWave<=-135;CosWave<=-375; end
    112:begin SinWave<=-147;CosWave<=-371; end
    113:begin SinWave<=-158;CosWave<=-366; end
    114:begin SinWave<=-170;CosWave<=-361; end
    115:begin SinWave<=-181;CosWave<=-356; end
    116:begin SinWave<=-192;CosWave<=-350; end
    117:begin SinWave<=-203;CosWave<=-343; end
    118:begin SinWave<=-214;CosWave<=-337; end
    119:begin SinWave<=-224;CosWave<=-330; end
    120:begin SinWave<=-235;CosWave<=-323; end
    121:begin SinWave<=-245;CosWave<=-315; end
    122:begin SinWave<=-254;CosWave<=-307; end
    123:begin SinWave<=-264;CosWave<=-299; end
    124:begin SinWave<=-273;CosWave<=-291; end
    125:begin SinWave<=-282;CosWave<=-282; end
    126:begin SinWave<=-291;CosWave<=-273; end
    127:begin SinWave<=-299;CosWave<=-264; end
    128:begin SinWave<=-307;CosWave<=-254; end
    129:begin SinWave<=-315;CosWave<=-245; end
    130:begin SinWave<=-323;CosWave<=-235; end
    131:begin SinWave<=-330;CosWave<=-224; end
    132:begin SinWave<=-337;CosWave<=-214; end
    133:begin SinWave<=-343;CosWave<=-203; end
    134:begin SinWave<=-350;CosWave<=-192; end
    135:begin SinWave<=-356;CosWave<=-181; end
    136:begin SinWave<=-361;CosWave<=-170; end
    137:begin SinWave<=-366;CosWave<=-158; end
    138:begin SinWave<=-371;CosWave<=-147; end
    139:begin SinWave<=-375;CosWave<=-135; end
    140:begin SinWave<=-379;CosWave<=-123; end
    141:begin SinWave<=-383;CosWave<=-111; end
    142:begin SinWave<=-386;CosWave<=-99; end
    143:begin SinWave<=-389;CosWave<=-87; end
    144:begin SinWave<=-392;CosWave<=-75; end
    145:begin SinWave<=-394;CosWave<=-62; end
    146:begin SinWave<=-396;CosWave<=-50; end
    147:begin SinWave<=-397;CosWave<=-38; end
    148:begin SinWave<=-398;CosWave<=-25; end
    149:begin SinWave<=-399;CosWave<=-13; end
    150:begin SinWave<=-399;CosWave<=0; end
    151:begin SinWave<=-399;CosWave<=13; end
    152:begin SinWave<=-398;CosWave<=25; end
    153:begin SinWave<=-397;CosWave<=38; end
    154:begin SinWave<=-396;CosWave<=50; end
    155:begin SinWave<=-394;CosWave<=62; end
    156:begin SinWave<=-392;CosWave<=75; end
    157:begin SinWave<=-389;CosWave<=87; end
    158:begin SinWave<=-386;CosWave<=99; end
    159:begin SinWave<=-383;CosWave<=111; end
    160:begin SinWave<=-379;CosWave<=123; end
    161:begin SinWave<=-375;CosWave<=135; end
    162:begin SinWave<=-371;CosWave<=147; end
    163:begin SinWave<=-366;CosWave<=158; end
    164:begin SinWave<=-361;CosWave<=170; end
    165:begin SinWave<=-356;CosWave<=181; end
    166:begin SinWave<=-350;CosWave<=192; end
    167:begin SinWave<=-343;CosWave<=203; end
    168:begin SinWave<=-337;CosWave<=214; end
    169:begin SinWave<=-330;CosWave<=224; end
    170:begin SinWave<=-323;CosWave<=235; end
    171:begin SinWave<=-315;CosWave<=245; end
    172:begin SinWave<=-307;CosWave<=254; end
    173:begin SinWave<=-299;CosWave<=264; end
    174:begin SinWave<=-291;CosWave<=273; end
    175:begin SinWave<=-282;CosWave<=282; end
    176:begin SinWave<=-273;CosWave<=291; end
    177:begin SinWave<=-264;CosWave<=299; end
    178:begin SinWave<=-254;CosWave<=307; end
    179:begin SinWave<=-245;CosWave<=315; end
    180:begin SinWave<=-235;CosWave<=323; end
    181:begin SinWave<=-224;CosWave<=330; end
    182:begin SinWave<=-214;CosWave<=337; end
    183:begin SinWave<=-203;CosWave<=343; end
    184:begin SinWave<=-192;CosWave<=350; end
    185:begin SinWave<=-181;CosWave<=356; end
    186:begin SinWave<=-170;CosWave<=361; end
    187:begin SinWave<=-158;CosWave<=366; end
    188:begin SinWave<=-147;CosWave<=371; end
    189:begin SinWave<=-135;CosWave<=375; end
    190:begin SinWave<=-123;CosWave<=379; end
    191:begin SinWave<=-111;CosWave<=383; end
    192:begin SinWave<=-99;CosWave<=386; end
    193:begin SinWave<=-87;CosWave<=389; end
    194:begin SinWave<=-75;CosWave<=392; end
    195:begin SinWave<=-62;CosWave<=394; end
    196:begin SinWave<=-50;CosWave<=396; end
    197:begin SinWave<=-38;CosWave<=397; end
    198:begin SinWave<=-25;CosWave<=398; end
    199:begin SinWave<=-13;CosWave<=399; end

    endcase
  end
endmodule // CarryWaveGen
